package router_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"   // Always first

  // ============================================================
  // 1. Configurations
  // ============================================================
  `include "src_agent_config.sv"
  `include "dst_agent_config.sv"
  `include "router_env_config.sv"

  // ============================================================
  // 2. Transaction classes
  // ============================================================
  `include "src_xtn.sv"
  `include "dst_xtn.sv"

  // ============================================================
  // 3. Sequences
  // ============================================================
  `include "src_seqs.sv"
  `include "dst_seqs.sv"

  // ============================================================
  // 4. Sequencers
  // ============================================================
  `include "src_seqr.sv"
  `include "dst_seqr.sv"

  // ============================================================
  // 5. Drivers
  // ============================================================
  `include "src_driver.sv"
  `include "dst_driver.sv"

  // ============================================================
  // 6. Monitors
  // ============================================================
  `include "src_mon.sv"
  `include "dst_mon.sv"

  // ============================================================
  // 7. Agents
  // ============================================================
  `include "src_agent.sv"
  `include "dst_agent.sv"

  // ============================================================
  // 8. Agent Tops
  // ============================================================


  // ============================================================
  // 9. Virtual Sequencer + Virtual Sequences
  // ============================================================
  `include "router_virtual_sequencer.sv"
	`include "src_agent_top.sv"
  `include "dst_agent_top.sv"
  `include "router_scoreboard.sv"

  // ============================================================
  // 10. Environment
  // ============================================================

 `include "router_virtual_sequence.sv"
  `include "router_env.sv"

  // ============================================================
  // 11. Test
  // ============================================================
  `include "router_test_lib.sv"

endpackage
